`ifndef MEMORY_V
`define MEMORY_V

module memory();

endmodule

`endif